--/////////////////////////////////////////////////////////////////////////////////////////
-- Company: University at Buffalo
-- Engineer: Thomas Mehok
-- 
-- Create Date:    11/26/2024
-- Module Name:    SPI_Snake_EE478Final
-- Project Name:   SPI_Snake_EE478Final 
-- Target Devices: ZYBO Z7
-- Tool versions:  ISE 14.1
-- Description: This is a demo for the Digilent PmodACL.  The SW inputs are
--					 used to select either the x-axis, y-axis, or z-axis data for
--					 display, and RST is used to reset the demo.
--
--					 There are four main components in this module, SPIcomponent, sel_Data,
--					 ClkDiv_5Hz, and ssdCtrl.  A START signal is generated by the ClkDiv_5Hz
--					 component, this signal is used to initiate a data transfer between the
--					 PmodACL and the Nexys3.

--					THOMAS NOTES: Unsure of what the 5Hz clock does in the grand sceme. From this main module it is sent into SPImaster
--								  It seems to. DOUBLE CHECK *************** it seems like it is reading the doing a reading at the 5hz speed.
--								  I do not know where this number is coming from 
--
--					 SPIcomponent receives the START signal, configures the PmodACL, and then
--					 receives data pertaining to all three axes.  The data is made available
--					 to the rest of the design on the xAxis, yAxis, and zAxis outputs.

--					THOMAS NOTES: At this point in the module It is confirmed that the start signal starts off our SPIMaster state machine.
--								  We may not need most parts of the module as the outputs or SPIcomponent give us the X-axis, Y-axis, and Z-axis data
--
--					 These outputs are then sent into the sel_Data component with the the status
--					 of switches SW1 and SW0 on the Nexys3. Depending on the configuration of
--					 these switches, one of the axes data will be selected for display on the
--					 seven segment display. The selected data is converted from 2's compliment
--					 to magnitude, and is then sent to the ssdCtrl where it is converted to a "g"
--					 value and displayed on the SSD with hundredths precision.
--
--					THOMAS NOTES: I will not need the sel_Data and the ssdCtrl module. They are for displaying the gravity value. It might be useful
--								  to looking these files in order to better understand their conversion. We may still need them to convert to the correct 
--								  a comparable value that will allow us to compare which axis has the most acceleration connected to it.
--
--					 To select an axis for display configure SW1 and SW0 on the Nexys3 as
--					 shown below.  LED LD0 will illuminate when the x-axis is selected,
--					 LD1 for y-aixs, and LD2 for z-axis.
--
--							SW1	SW0	|	SSD Output	|	LD2	|	LD1	|	LD0
--							------------------------------------------------------
--							off	off	|	x-axis		|	off	|	off	|	on
--							off	on	|	y-axis		|	off	|	on	|	off
--							on	on	|	x-axis		|	off	|	off	|	on
--							on	off	|	z-axis		|	on	|	off	|	off

--					THOMAS NOTES: Good chance we will not use these buttons as all but still we wan to convert these numbers.

--					THOMAS NOTES: We are going to need to add in more modules of our own in order to output the values our partner is looking for 
--								  the video game


-- ================================================================================================================================
--											DOMINANT DIRECTION MODULE
-- ================================================================================================================================
--					The DDmodule will allow us to get the most dominant of the current axis in terms of acceleration with a small buffer 
--					in order to not be fragile to any movment when trying to control the snake. This buffer will act as almost debouncing
--					

--  Inputs:
--		CLK				Onboard system clock
--		RST				Resets the demo
--		SW<0>				Selects y-axis data for display
--		SW<1>				Selects z-axis data for display
--		SDI				Serial Data In
--
--  Outputs:
--		SDO				Serial Data Out
--		SCLK				Serial Clock
--		SS					Slave Select

--		THOMAS NOTES: I do not believe this output will be nessasary******************
--		AN				Anodes on SSD
--		SEG				Cathodes on SSD
--		DOT				Cathode for decimal on SSD

--		THOMAS NOTES: This is going to be the LED we output to the ZYBO board to all the user to confirm what direction they are going
--		LED				LEDs on ZYBO Z7
--
-- Revision History: 
-- 						Revision 0.01 - File Created (Josh Sackos)
--/////////////////////////////////////////////////////////////////////////////////////////
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.std_logic_arith.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- ====================================================================================
-- 										  Define Module
-- ====================================================================================
entity PmodACL_Demo is
    Port ( 
		   CLK : in  STD_LOGIC;
           RST : in  STD_LOGIC;
           --SW : in  STD_LOGIC_VECTOR (1 downto 0);
           SDI : in  STD_LOGIC;
           SDO : out  STD_LOGIC;
           SCLK : out  STD_LOGIC;
           SS : out  STD_LOGIC;
		   --LEDout : out STD_LOGIC_VECTOR(3 downto 0);
           --AN : out  STD_LOGIC_VECTOR (3 downto 0);
           --SEG : out  STD_LOGIC_VECTOR (6 downto 0);
           --DOT : out  STD_LOGIC;
           LED : out  STD_LOGIC_VECTOR (3 downto 0)
		   );
end PmodACL_Demo;

architecture Behavioral of PmodACL_Demo is


--  ===================================================================================
-- 							  				  Components
--  ===================================================================================

		-- **********************************************
		-- 		 			 Select Data
		--					Will not need
		-- **********************************************
		-- component sel_Data Port(
		-- 			CLK : in  STD_LOGIC;
		-- 			RST : in  STD_LOGIC;
		-- 			SW : in STD_LOGIC_VECTOR(1 downto 0);
		-- 			xAxis : in  STD_LOGIC_VECTOR (9 downto 0);
		-- 			yAxis : in  STD_LOGIC_VECTOR (9 downto 0);
		-- 			zAxis : in  STD_LOGIC_VECTOR (9 downto 0);
		-- 			DOUT : out  STD_LOGIC_VECTOR (9 downto 0);
		-- 			LED : out  STD_LOGIC_VECTOR (2 downto 0)
		-- );
		-- end component;

		-- **********************************************
		-- 		 Seven Segment Display Controller
		-- **********************************************
		component SPIcomponent
			Port ( CLK : in  STD_LOGIC;
					 RST : in  STD_LOGIC;
					 START : in STD_LOGIC;
					 SDI : in  STD_LOGIC;
					 SDO : out  STD_LOGIC;
					 SCLK : out  STD_LOGIC;
					 SS : out  STD_LOGIC;
					 xAxis : out STD_LOGIC_VECTOR(9 downto 0);
					 yAxis : out STD_LOGIC_VECTOR(9 downto 0);
					 zAxis : out STD_LOGIC_VECTOR(9 downto 0)
			 );
		end component;

		-- **********************************************
		-- 		 Seven Segment Display Controller
		--			Will not need this module 
		-- **********************************************
		-- component ssdCtrl
		-- 	 Port ( CLK : in  STD_LOGIC;
		-- 			  RST : in  STD_LOGIC;
		-- 			  DIN : in  STD_LOGIC_VECTOR (9 downto 0);
		-- 			  AN : out  STD_LOGIC_VECTOR (3 downto 0);
		-- 			  SEG : out  STD_LOGIC_VECTOR (6 downto 0);
		-- 			  DOT : out STD_LOGIC
		-- 	 );
		-- end component;

		-- **********************************************
		-- 				5Hz Clock Divider
		-- **********************************************
		component ClkDiv_5Hz
			Port (  
					CLK : in  STD_LOGIC;
					RST : in STD_LOGIC;
					CLKOUT : inout STD_LOGIC
				);
		end component;

		-- **********************************************
		--				DOMINANT DIRECTION MODULE
		-- **********************************************

		component DDmodule
			Port (
					CLK : 		in STD_LOGIC;
					DDirection: out STD_LOGIC_VECTOR(3 downto 0);
					xAxis : 	in STD_LOGIC_VECTOR(9 downto 0);
					yAxis :		in STD_LOGIC_VECTOR(9 downto 0);
					zAxis : 	in STD_LOGIC_VECTOR(9 downto 0)
			);
		end component;

-- ====================================================================================
-- 							       Signals and Constants
-- ====================================================================================

		signal xAxis : STD_LOGIC_VECTOR(9 downto 0);		-- x-axis data from PmodACL
		signal yAxis : STD_LOGIC_VECTOR(9 downto 0);		-- y-axis data from PmodACL
		signal zAxis : STD_LOGIC_VECTOR(9 downto 0);		-- z-axis data from PmodACL

		signal selData : STD_LOGIC_VECTOR(9 downto 0);	-- Data selected to display

		signal START : STD_LOGIC;								-- Data Transfer Request Signal

-- ////////////////////////////////////////////////////////////////////////////////////////////////////////
--											Start of Thomas Mehok Signals
-- ////////////////////////////////////////////////////////////////////////////////////////////////////////
		--signal LEDout : STD_LOGIC_VECTOR(3 downto 0);		-- This signal represents what LED will be lit up on the board itself

--  ===================================================================================
-- 							  				Implementation
--  ===================================================================================
begin

			-------------------------------------------------
			--	Select Display Data and Convert to Magnitude
			-------------------------------------------------
			-- SDATA : sel_Data port map(
			-- 				CLK=>CLK,
			-- 				RST=>RST,
			-- 				SW=>SW,
			-- 				xAxis=>xAxis,
			-- 				yAxis=>yAxis,
			-- 				zAxis=>zAxis,
			-- 				DOUT=>selData,
			-- 				LED=>LED
			-- );

			-------------------------------------------------
			--		 			 Interfaces PmodACL
			-------------------------------------------------
			SPI : SPIcomponent port map(
							CLK=>CLK,
							RST=>RST,
							START=>START,
							SDI=>SDI,
							SDO=>SDO,
							SCLK=>SCLK,
							SS=>SS,
							xAxis=>xAxis,
							yAxis=>yAxis,
							zAxis=>zAxis
			);

			-------------------------------------------------
			--		 	 Formats Data and Displays on SSD
			-------------------------------------------------
			-- Disp : ssdCtrl port map(
			-- 				CLK=>CLK,
			-- 				RST=>RST,
			-- 				DIN=>selData(9 downto 0),
			-- 				AN=>AN,
			-- 				SEG=>SEG,
			-- 				DOT=>DOT
			-- );

			-------------------------------------------------
			--	 Generates a 5Hz Data Transfer Request Signal
			-------------------------------------------------
			genStart : ClkDiv_5Hz port map(
							CLK=>CLK,
							RST=>RST,
							CLKOUT=>START
			);

			LED_DOM : DDmodule port map (
					CLK => CLK,
					DDirection => LED,
					xAxis => xAxis,
					yAxis => yAxis,
					zAxis => zAxis
			);

end Behavioral;

